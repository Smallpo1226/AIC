
.SUBCKT Diff_AMP VDD VSS Vb Vin Vip Voutn Voutp
CC1 Voutn VSS 1p 
CC0 Voutp VSS 1p 
RR1 VDD Voutp 100.690K
RR0 VDD Voutn 100.690K
MM3 net26 Vb VSS VSS N_18 W=5.166u  L=3u m=35
MM2 Voutp Vin net26 VSS N_18 W=14.685u  L=4.4u m=8
MM1 Voutn Vip net26 VSS N_18 W=14.685u  L=4.4u m=8
.ENDS

